library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- First entity
entity decimal_to_sseg is
    port (dec_in   : in  std_logic_vector(3 downto 0);  
			 sseg_out : out std_logic_vector(0 to 6));
end entity decimal_to_sseg;

architecture behaviour of decimal_to_sseg is
begin
	with dec_in select
		sseg_out <= "0000001" when "0000",
					   "1001111" when "0001",
						"0010010" when "0010",
						"0000110" when "0011",
						"1001100" when "0100",
						"0100100" when "0101",
						"0100000" when "0110",
						"0001111" when "0111",
						"0000000" when "1000",
						"0000100" when "1001",
						"1111111" when others;
end behaviour;